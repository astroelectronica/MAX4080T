.title KiCad schematic
.include "C:/AE/MAX4080T/_models/C2012C0G2E102J085AA_p.mod"
.include "C:/AE/MAX4080T/_models/C2012X7R2A104K125AA_p.mod"
.include "C:/AE/MAX4080T/_models/C2012X7R2E103K125AA_p.mod"
.include "C:/AE/MAX4080T/_models/C3216X5R1H106M160AB_p.mod"
.include "C:/AE/MAX4080T/_models/MAX4080T.FAM"
R1 /VOUT /VIN {RSNS}
V1 /VIN 0 {VSOURCE}
XU1 /VIN 0 C3216X5R1H106M160AB_p
XU2 /VIN 0 C2012X7R2A104K125AA_p
I1 /VOUT 0 {ILOAD}
XU4 /RSP /VIN unconnected-_U4-NC-Pad3_ 0 /VOCM unconnected-_U4-NC-Pad6_ unconnected-_U4-NC-Pad7_ /RSN MAX4080T
R5 /VOCM /OUT {RLPF}
R4 /VOUT /RSN {RLIM}
R3 /VIN /RSP {RLIM}
R2 /VOUT /VIN {RSNS}
XU3 /RSN /RSP C2012C0G2E102J085AA_p
XU5 0 /OUT C2012X7R2E103K125AA_p
.end
